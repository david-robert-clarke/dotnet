-- Final Year Project
-- By David.R.Clarke
-- Created on 10_12_2000
-- Updated on 11_12_2000
Library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
--
ENTITY Answer_Store IS
--PORT (D : IN STD_LOGIC, CLK : IN STD_LOGIC; Q : OUT STD_LOGIC_VECTOR (19 DOWNTO 0));
PORT (CE,CLR          : IN STD_LOGIC;
      SOP_IN          : IN STD_LOGIC_VECTOR (4 downto 0); 
      LATCH_MEM       : IN STD_LOGIC_VECTOR (3 downto 0); 
      A0B0_A1B2, A0B1_A1B3, A2B0_A3B2, A2B1_A3B3 : OUT STD_LOGIC_VECTOR (4 downto 0));
END ENTITY Answer_Store;
--
ARCHITECTURE STRUCTURAL OF Answer_Store IS

COMPONENT FDCE IS
Port (D, C, CLR, CE : IN STD_LOGIC; Q : OUT STD_LOGIC);
END COMPONENT FDCE;

-- SIGNAL SOP_BUS_IN : STD_LOGIC_VECTOR (4 downto 0); 
--       LATCH_BUS  : STD_LOGIC_VECTOR (3 downto 0); 
--       ANS_BUS_3, ANS_BUS_2, ANS_BUS_1, ANS_BUS_0 : STD_LOGIC_VECTOR (4 downto 0));

BEGIN

FDCE19 : FDCE PORT MAP (D => SOP_IN(4), C => LATCH_MEM(3), Q => A0B0_A1B2(4), CLR => CLR, CE => CE);
FDCE18 : FDCE PORT MAP (D => SOP_IN(3), C => LATCH_MEM(3), Q => A0B0_A1B2(3), CLR => CLR, CE => CE);
FDCE17 : FDCE PORT MAP (D => SOP_IN(2), C => LATCH_MEM(3), Q => A0B0_A1B2(2), CLR => CLR, CE => CE);
FDCE16 : FDCE PORT MAP (D => SOP_IN(1), C => LATCH_MEM(3), Q => A0B0_A1B2(1), CLR => CLR, CE => CE);
FDCE15 : FDCE PORT MAP (D => SOP_IN(0), C => LATCH_MEM(3), Q => A0B0_A1B2(0), CLR => CLR, CE => CE);
FDCE14 : FDCE PORT MAP (D => SOP_IN(4), C => LATCH_MEM(2), Q => A0B1_A1B3(4), CLR => CLR, CE => CE);
FDCE13 : FDCE PORT MAP (D => SOP_IN(3), C => LATCH_MEM(2), Q => A0B1_A1B3(3), CLR => CLR, CE => CE);
FDCE12 : FDCE PORT MAP (D => SOP_IN(2), C => LATCH_MEM(2), Q => A0B1_A1B3(2), CLR => CLR, CE => CE);
FDCE11 : FDCE PORT MAP (D => SOP_IN(1), C => LATCH_MEM(2), Q => A0B1_A1B3(1), CLR => CLR, CE => CE);
FDCE10 : FDCE PORT MAP (D => SOP_IN(0), C => LATCH_MEM(2), Q => A0B1_A1B3(0), CLR => CLR, CE => CE);
FDCE9  : FDCE PORT MAP (D => SOP_IN(4), C => LATCH_MEM(1), Q => A2B0_A3B2(4), CLR => CLR, CE => CE);
FDCE8  : FDCE PORT MAP (D => SOP_IN(3), C => LATCH_MEM(1), Q => A2B0_A3B2(3), CLR => CLR, CE => CE);
FDCE7  : FDCE PORT MAP (D => SOP_IN(2), C => LATCH_MEM(1), Q => A2B0_A3B2(2), CLR => CLR, CE => CE);
FDCE6  : FDCE PORT MAP (D => SOP_IN(1), C => LATCH_MEM(1), Q => A2B0_A3B2(1), CLR => CLR, CE => CE);
FDCE5  : FDCE PORT MAP (D => SOP_IN(0), C => LATCH_MEM(1), Q => A2B0_A3B2(0), CLR => CLR, CE => CE);
FDCE4  : FDCE PORT MAP (D => SOP_IN(4), C => LATCH_MEM(0), Q => A2B1_A3B3(4), CLR => CLR, CE => CE);
FDCE3  : FDCE PORT MAP (D => SOP_IN(3), C => LATCH_MEM(0), Q => A2B1_A3B3(3), CLR => CLR, CE => CE);
FDCE2  : FDCE PORT MAP (D => SOP_IN(2), C => LATCH_MEM(0), Q => A2B1_A3B3(2), CLR => CLR, CE => CE);
FDCE1  : FDCE PORT MAP (D => SOP_IN(1), C => LATCH_MEM(0), Q => A2B1_A3B3(1), CLR => CLR, CE => CE);
FDCE0  : FDCE PORT MAP (D => SOP_IN(0), C => LATCH_MEM(0), Q => A2B1_A3B3(0), CLR => CLR, CE => CE);

END ARCHITECTURE STRUCTURAL;

 

-- Created by David Clarke for the RS232 assignment
library IEEE;
use IEEE.std_logic_1164.all;

entity OR5 is
    port (a : in STD_LOGIC; b : in STD_LOGIC; c: in STD_LOGIC; 
          d : in STD_LOGIC; e : in STD_LOGIC; z: out STD_LOGIC);
end OR5;

architecture behavioural of OR5 is
begin
  
  z <= a or b or c or d or e;
  
end behavioural;

-- Final Year project messaround
-- Created by David Clarke
Library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE WORK.MATRIX_PACKAGE.ALL;

ENTITY MUL_2BIT IS 
	PORT (A, B : IN U_TWO_BITS; Z : OUT NIBBLE);
END ENTITY MUL_2BIT;
--
ARCHITECTURE BEHAVIOURAL OF MUL_2BIT IS
BEGIN

	Z  <= CONV_STD_LOGIC_VECTOR((A*B), 4);

END ARCHITECTURE BEHAVIOURAL;

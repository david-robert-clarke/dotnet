-- ACTIVE-CAD-2-VHDL, 2.5.5.67, Wed Nov 15 18:47:52 2000

library IEEE;
use IEEE.std_logic_1164.all;

entity wholesystem is port (
	Q : out STD_LOGIC_VECTOR (15 downto 0);
	X36_NET00043_X95 : out STD_LOGIC;
	X36_NET00044_X95 : out STD_LOGIC;
	X36_NET00052_X95 : out STD_LOGIC;
	X36_NET00053_X95 : in STD_LOGIC;
	X36_NET00054_X95 : out STD_LOGIC;
	X36_NET00055_X95 : in STD_LOGIC;
	X36_NET00056_X95 : in STD_LOGIC;
	X36_NET00058_X95 : out STD_LOGIC
); end WHOLESYSTEM;

architecture SCHEMATIC of WHOLESYSTEM is

--COMPONENTS

component CONTROLBEAST port (
	CLK : in STD_LOGIC;
	CLR : in STD_LOGIC;
	PTEN : out STD_LOGIC;
	UP : out STD_LOGIC;
	CDDEN : out STD_LOGIC;
	CT1EN : out STD_LOGIC;
	DECEN : out STD_LOGIC;
	LOAD : out STD_LOGIC;
	CT1Z : in STD_LOGIC;
	S : in STD_LOGIC
); end component;

component CB16CLED port (
	D : in STD_LOGIC_VECTOR (15 downto 0);
	Q : out STD_LOGIC_VECTOR (15 downto 0);
	C : in STD_LOGIC;
	CE : in STD_LOGIC;
	CEO : out STD_LOGIC;
	CLR : in STD_LOGIC;
	L : in STD_LOGIC;
	TC : out STD_LOGIC;
	UP : in STD_LOGIC
); end component;

component DECODER port (
	B6 : in STD_LOGIC;
	B7 : in STD_LOGIC;
	B10 : in STD_LOGIC;
	B8 : in STD_LOGIC;
	B9 : in STD_LOGIC;
	B11 : in STD_LOGIC;
	DECEN : in STD_LOGIC;
	S300 : out STD_LOGIC;
	S2400 : out STD_LOGIC;
	S4800 : out STD_LOGIC;
	S600 : out STD_LOGIC;
	S1200 : out STD_LOGIC;
	S9600 : out STD_LOGIC;
	S19200 : out STD_LOGIC;
	RESET : in STD_LOGIC
); end component;

component CDDECODE port (
	CNT : out STD_LOGIC_VECTOR (15 downto 0);
	CDDEN : in STD_LOGIC;
	RESET : in STD_LOGIC;
	S19200 : in STD_LOGIC;
	S4800 : in STD_LOGIC;
	S9600 : in STD_LOGIC;
	S600 : in STD_LOGIC;
	S2400 : in STD_LOGIC;
	S1200 : in STD_LOGIC;
	S300 : in STD_LOGIC
); end component;

component PARITY_TEST port (
	EVEN : out STD_LOGIC;
	ODD : out STD_LOGIC;
	PTEN : in STD_LOGIC;
	RESET : in STD_LOGIC;
	S : in STD_LOGIC
); end component;

component OBUF port (
	I : in STD_LOGIC;
	O : out STD_LOGIC
); end component;

component IBUF port (
	I : in STD_LOGIC;
	O : out STD_LOGIC
); end component;

component PINOUTDECODE port (
	RESET : in STD_LOGIC;
	S19200 : in STD_LOGIC;
	S4800 : in STD_LOGIC;
	S9600 : in STD_LOGIC;
	S2400 : in STD_LOGIC;
	S1200 : in STD_LOGIC;
	S600 : in STD_LOGIC;
	S300 : in STD_LOGIC;
	S6 : out STD_LOGIC;
	S4 : out STD_LOGIC;
	S5 : out STD_LOGIC
); end component;

component INV port (
	I : in STD_LOGIC;
	O : out STD_LOGIC
); end component;

--SIGNALS

signal X36_NET00033_X95 : STD_LOGIC;
signal X36_NET00034_X95 : STD_LOGIC;
signal X36_NET00035_X95 : STD_LOGIC;
signal S : STD_LOGIC;
signal X36_NET00037_X95 : STD_LOGIC;
signal X36_NET00038_X95 : STD_LOGIC;
signal X36_NET00039_X95 : STD_LOGIC;
signal X36_NET00040_X95 : STD_LOGIC;
signal X36_NET00041_X95 : STD_LOGIC;
signal X36_NET00042_X95 : STD_LOGIC;
signal X36_NET00045_X95 : STD_LOGIC;
signal X36_NET00046_X95 : STD_LOGIC;
signal X36_NET00047_X95 : STD_LOGIC;
signal X36_NET00048_X95 : STD_LOGIC;
signal X36_NET00049_X95 : STD_LOGIC;
signal X36_NET00050_X95 : STD_LOGIC;
signal X36_NET00051_X95 : STD_LOGIC;
signal X36_NET00057_X95 : STD_LOGIC;
signal X36_NET00059_X95 : STD_LOGIC;
signal X36_NET00060_X95 : STD_LOGIC;
signal X36_NET00061_X95 : STD_LOGIC;
signal X36_NET00062_X95 : STD_LOGIC;
signal X36_NET00063_X95 : STD_LOGIC;
signal Q11_ASSIGN_B11 : STD_LOGIC;
signal Q10_ASSIGN_B10 : STD_LOGIC;
signal Q9_ASSIGN_B9 : STD_LOGIC;
signal Q8_ASSIGN_B8 : STD_LOGIC;
signal Q7_ASSIGN_B7 : STD_LOGIC;
signal Q6_ASSIGN_B6 : STD_LOGIC;
signal X36_NET00043_ASSIGN_OPAD : STD_LOGIC;
signal X36_NET00044_ASSIGN_OPAD : STD_LOGIC;
signal X36_NET00052_ASSIGN_OPAD : STD_LOGIC;
signal X36_NET00053_ASSIGN_IPAD : STD_LOGIC;
signal X36_NET00054_ASSIGN_OPAD : STD_LOGIC;
signal X36_NET00055_ASSIGN_IPAD : STD_LOGIC;
signal X36_NET00056_ASSIGN_IPAD : STD_LOGIC;
signal X36_NET00058_ASSIGN_OPAD : STD_LOGIC;
signal X36_I31_GTS_I : STD_LOGIC;
signal X36_I33_GTS_I : STD_LOGIC;
signal X36_I32_GTS_I : STD_LOGIC;
signal X36_I26_GTS_I : STD_LOGIC;
signal X36_I25_GTS_I : STD_LOGIC;

signal CNT : STD_LOGIC_VECTOR (15 downto 0);

--ATRIBUTES





begin

--SIGNAL ASSIGNMENTS

Q(11) <= Q11_ASSIGN_B11;
Q(10) <= Q10_ASSIGN_B10;
Q(9) <= Q9_ASSIGN_B9;
Q(8) <= Q8_ASSIGN_B8;
Q(7) <= Q7_ASSIGN_B7;
Q(6) <= Q6_ASSIGN_B6;
X36_NET00043_X95 <= X36_NET00043_ASSIGN_OPAD;
X36_NET00044_X95 <= X36_NET00044_ASSIGN_OPAD;
X36_NET00052_X95 <= X36_NET00052_ASSIGN_OPAD;
X36_NET00053_ASSIGN_IPAD <= X36_NET00053_X95;
X36_NET00054_X95 <= X36_NET00054_ASSIGN_OPAD;
X36_NET00055_ASSIGN_IPAD <= X36_NET00055_X95;
X36_NET00056_ASSIGN_IPAD <= X36_NET00056_X95;
X36_NET00058_X95 <= X36_NET00058_ASSIGN_OPAD;

--COMPONENT INSTANCES

H1 : CONTROLBEAST port map(
	CLK => X36_NET00037_X95,
	CLR => X36_NET00035_X95,
	PTEN => X36_NET00033_X95,
	UP => X36_NET00040_X95,
	CDDEN => X36_NET00039_X95,
	CT1EN => X36_NET00042_X95,
	DECEN => X36_NET00063_X95,
	LOAD => X36_NET00041_X95,
	CT1Z => X36_NET00038_X95,
	S => S
);
X36_I1 : CB16CLED port map(
	D(15) => CNT(15),
	D(14) => CNT(14),
	D(13) => CNT(13),
	D(12) => CNT(12),
	D(11) => CNT(11),
	D(10) => CNT(10),
	D(9) => CNT(9),
	D(8) => CNT(8),
	D(7) => CNT(7),
	D(6) => CNT(6),
	D(5) => CNT(5),
	D(4) => CNT(4),
	D(3) => CNT(3),
	D(2) => CNT(2),
	D(1) => CNT(1),
	D(0) => CNT(0),
	Q(15) => Q(15),
	Q(14) => Q(14),
	Q(13) => Q(13),
	Q(12) => Q(12),
	Q(11) => Q11_ASSIGN_B11,
	Q(10) => Q10_ASSIGN_B10,
	Q(9) => Q9_ASSIGN_B9,
	Q(8) => Q8_ASSIGN_B8,
	Q(7) => Q7_ASSIGN_B7,
	Q(6) => Q6_ASSIGN_B6,
	Q(5) => Q(5),
	Q(4) => Q(4),
	Q(3) => Q(3),
	Q(2) => Q(2),
	Q(1) => Q(1),
	Q(0) => Q(0),
	C => X36_NET00037_X95,
	CE => X36_NET00042_X95,
	CEO => X36_NET00038_X95,
	CLR => X36_NET00035_X95,
	L => X36_NET00041_X95,
	UP => X36_NET00040_X95
);
U1 : DECODER port map(
	B6 => Q6_ASSIGN_B6,
	B7 => Q7_ASSIGN_B7,
	B10 => Q10_ASSIGN_B10,
	B8 => Q8_ASSIGN_B8,
	B9 => Q9_ASSIGN_B9,
	B11 => Q11_ASSIGN_B11,
	DECEN => X36_NET00063_X95,
	S300 => X36_NET00045_X95,
	S2400 => X36_NET00048_X95,
	S4800 => X36_NET00049_X95,
	S600 => X36_NET00046_X95,
	S1200 => X36_NET00047_X95,
	S9600 => X36_NET00050_X95,
	S19200 => X36_NET00051_X95,
	RESET => X36_NET00035_X95
);
U2 : CDDECODE port map(
	CNT(15) => CNT(15),
	CNT(14) => CNT(14),
	CNT(13) => CNT(13),
	CNT(12) => CNT(12),
	CNT(11) => CNT(11),
	CNT(10) => CNT(10),
	CNT(9) => CNT(9),
	CNT(8) => CNT(8),
	CNT(7) => CNT(7),
	CNT(6) => CNT(6),
	CNT(5) => CNT(5),
	CNT(4) => CNT(4),
	CNT(3) => CNT(3),
	CNT(2) => CNT(2),
	CNT(1) => CNT(1),
	CNT(0) => CNT(0),
	CDDEN => X36_NET00039_X95,
	RESET => X36_NET00035_X95,
	S19200 => X36_NET00051_X95,
	S4800 => X36_NET00049_X95,
	S9600 => X36_NET00050_X95,
	S600 => X36_NET00046_X95,
	S2400 => X36_NET00048_X95,
	S1200 => X36_NET00047_X95,
	S300 => X36_NET00045_X95
);
U3 : PARITY_TEST port map(
	EVEN => X36_NET00062_X95,
	ODD => X36_NET00034_X95,
	PTEN => X36_NET00033_X95,
	RESET => X36_NET00035_X95,
	S => S
);
X36_I31 : OBUF port map(
	I => X36_NET00060_X95,
	O => X36_NET00044_ASSIGN_OPAD
);
X36_I33 : OBUF port map(
	I => X36_NET00061_X95,
	O => X36_NET00043_ASSIGN_OPAD
);
X36_I32 : OBUF port map(
	I => X36_NET00059_X95,
	O => X36_NET00052_ASSIGN_OPAD
);
X36_I26 : OBUF port map(
	I => X36_NET00062_X95,
	O => X36_NET00054_ASSIGN_OPAD
);
X36_I24 : IBUF port map(
	I => X36_NET00055_ASSIGN_IPAD,
	O => X36_NET00035_X95
);
U4 : PINOUTDECODE port map(
	RESET => X36_NET00035_X95,
	S19200 => X36_NET00051_X95,
	S4800 => X36_NET00049_X95,
	S9600 => X36_NET00050_X95,
	S2400 => X36_NET00048_X95,
	S1200 => X36_NET00047_X95,
	S600 => X36_NET00046_X95,
	S300 => X36_NET00045_X95,
	S6 => X36_NET00059_X95,
	S4 => X36_NET00061_X95,
	S5 => X36_NET00060_X95
);
X36_I23 : IBUF port map(
	I => X36_NET00056_ASSIGN_IPAD,
	O => X36_NET00057_X95
);
X36_I19 : IBUF port map(
	I => X36_NET00053_ASSIGN_IPAD,
	O => X36_NET00037_X95
);
X36_I25 : OBUF port map(
	I => X36_NET00034_X95,
	O => X36_NET00058_ASSIGN_OPAD
);
X36_I35 : INV port map(
	I => X36_NET00057_X95,
	O => S
);

end SCHEMATIC;


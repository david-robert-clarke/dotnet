-- Final Year project 
-- By David Clarke
-- Created 30_1_2001
Library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE WORK.MATRIX_PACKAGE.ALL;

ENTITY MUL_TWO_BITS IS 
	PORT (A, B : IN U_TWO_BITS; Z : OUT NIBBLE);
END ENTITY MUL_TWO_BITS;
--
ARCHITECTURE BEHAVIOURAL OF MUL_TWO_BITS IS
BEGIN

	Z  <= CONV_STD_LOGIC_VECTOR((A*B), 4);
	
END ARCHITECTURE BEHAVIOURAL;

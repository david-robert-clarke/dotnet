-- Created by David Clarke for the RS232 assignment
library IEEE;
use IEEE.std_logic_1164.all;

entity OR2 is
    port (a: in STD_LOGIC; b: in STD_LOGIC;
          z: out STD_LOGIC);
end OR2;

architecture behavioural of OR2 is
begin
  
  z <= a or b;
  
end behavioural;

-- Created by David Clarke for the RS232 assignment
library IEEE;
use IEEE.std_logic_1164.all;

entity M2_1B1 is port (
	D0 : in STD_LOGIC;
	D1 : in STD_LOGIC;
	O : out STD_LOGIC;
	S0 : in STD_LOGIC
); end M2_1B1;

architecture SCHEMATIC of M2_1B1 is

--COMPONENTS

component AND2B2 port (
	b : in STD_LOGIC;
	a : in STD_LOGIC;
	z : out STD_LOGIC
); end component;

component OR2 port (
	b : in STD_LOGIC;
	a : in STD_LOGIC;
	z : out STD_LOGIC
); end component;

component AND2 port (
	b : in STD_LOGIC;
	a : in STD_LOGIC;
	z : out STD_LOGIC
); end component;

--SIGNALS

signal M0 : STD_LOGIC;
signal M1 : STD_LOGIC;

--ATRIBUTES

begin

--SIGNAL ASSIGNMENTS


--COMPONENT INSTANCES

X36_1I7 : AND2B2 port map(
	b => S0,
	a => D0,
	z => M0
);
X36_1I8 : OR2 port map(
	b => M1,
	a => M0,
	z => O
);
X36_1I9 : AND2 port map(
	b => D1,
	a => S0,
	z => M1
);

end SCHEMATIC;

-- Created by David Clarke for the RS232 assignment
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

Entity AND2B1 IS
Port (a,b : IN std_logic; z : OUT std_logic);
End Entity AND2B1;

Architecture Behavioural OF AND2B1 IS
Begin
   z <= a AND (NOT b);
End Architecture Behavioural;

-- Final Year Project
-- By David Clarke
-- Created on 13_12_2000
-- Updated on 14_12_2000
library IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.std_logic_arith.ALL;

package MATRIX_PACKAGE IS
 subtype One_Bit           is STD_LOGIC;
 subtype Two_Bits          is STD_LOGIC_VECTOR (1 downto 0);
 subtype Three_Bits        is STD_LOGIC_VECTOR (2 downto 0);
 subtype NIBBLE            is STD_LOGIC_VECTOR (3 downto 0);
 subtype Five_Bits         is STD_LOGIC_VECTOR (4 downto 0);
 subtype Six_Bits          is STD_LOGIC_VECTOR (5 downto 0);
 subtype Seven_Bits        is STD_LOGIC_VECTOR (6 downto 0);
 subtype Byte              is STD_LOGIC_VECTOR (7 downto 0);
 subtype Nine_Bits         is STD_LOGIC_VECTOR (8 downto 0);
 subtype Ten_Bits          is STD_LOGIC_VECTOR (9 downto 0);
 subtype Eleven_Bits       is STD_LOGIC_VECTOR (10 downto 0);
 subtype Twelve_Bits       is STD_LOGIC_VECTOR (11 downto 0);
 subtype Thirteen_Bits     is STD_LOGIC_VECTOR (12 downto 0);
 subtype Fourteen_Bits     is STD_LOGIC_VECTOR (13 downto 0);
 subtype Fifteen_Bits      is STD_LOGIC_VECTOR (14 downto 0);
 subtype Word              is STD_LOGIC_VECTOR (15 downto 0);
 subtype Seventeen_Bits    is STD_LOGIC_VECTOR (16 downto 0);
 subtype Eigthteen_Bits    is STD_LOGIC_VECTOR (17 downto 0);
 subtype Nineteen_Bits     is STD_LOGIC_VECTOR (18 downto 0);
 subtype Twenty_Bits       is STD_LOGIC_VECTOR (19 downto 0);
 subtype Twenty1_Bits	   is STD_LOGIC_VECTOR (20 downto 0);
 subtype Twenty2_Bits      is STD_LOGIC_VECTOR (21 downto 0);
 subtype Twenty3_Bits      is STD_LOGIC_VECTOR (22 downto 0);
 subtype Twenty4_Bits      is STD_LOGIC_VECTOR (23 downto 0);
 subtype Twenty5_Bits      is STD_LOGIC_VECTOR (24 downto 0);
 subtype Twenty6_Bits      is STD_LOGIC_VECTOR (25 downto 0);
 subtype Twenty7_Bits      is STD_LOGIC_VECTOR (26 downto 0);
 subtype Twenty8_Bits      is STD_LOGIC_VECTOR (27 downto 0);
 subtype Twenty9_Bits      is STD_LOGIC_VECTOR (28 downto 0);
 subtype Thirty_Bits       is STD_LOGIC_VECTOR (29 downto 0);
 subtype Thirty1_Bits      is STD_LOGIC_VECTOR (30 downto 0);
 subtype Long_Word         is STD_LOGIC_VECTOR (31 downto 0);
 subtype Thirty3_Bits      is STD_LOGIC_VECTOR (32 downto 0);
 subtype Thirty4_Bits      is STD_LOGIC_VECTOR (33 downto 0);
 subtype Thirty5_Bits      is STD_LOGIC_VECTOR (34 downto 0);
 subtype Thirty6_Bits      is STD_LOGIC_VECTOR (35 downto 0);
 subtype Thirty7_Bits      is STD_LOGIC_VECTOR (36 downto 0);
 subtype Thirty8_Bits      is STD_LOGIC_VECTOR (37 downto 0);
 subtype Thirty9_Bits      is STD_LOGIC_VECTOR (38 downto 0);
 subtype Forty_Bits       is STD_LOGIC_VECTOR (39 downto 0);
 subtype Forty1_Bits      is STD_LOGIC_VECTOR (40 downto 0);
 subtype Forty2_Bits      is STD_LOGIC_VECTOR (41 downto 0);
 subtype Forty3_Bits      is STD_LOGIC_VECTOR (42 downto 0);
 subtype Forty4_Bits      is STD_LOGIC_VECTOR (43 downto 0);
 subtype Forty5_Bits      is STD_LOGIC_VECTOR (44 downto 0);
-- 
 subtype U_Two_Bits          is UNSIGNED (1 downto 0);
 subtype U_Three_Bits        is UNSIGNED (2 downto 0);
 subtype U_NIBBLE            is UNSIGNED (3 downto 0);
 subtype U_Five_Bits         is UNSIGNED (4 downto 0);
 subtype U_Six_Bits          is UNSIGNED (5 downto 0);
 subtype U_Seven_Bits        is UNSIGNED (6 downto 0);
 subtype U_Byte              is UNSIGNED (7 downto 0);
 subtype U_Nine_Bits         is UNSIGNED (8 downto 0);
 subtype U_Ten_Bits          is UNSIGNED (9 downto 0);
 subtype U_Eleven_Bits       is UNSIGNED (10 downto 0);
 subtype U_Twelve_Bits       is UNSIGNED (11 downto 0);
 subtype U_Thirteen_Bits     is UNSIGNED (12 downto 0);
 subtype U_Fourteen_Bits     is UNSIGNED (13 downto 0);
 subtype U_Fifteen_Bits      is UNSIGNED (14 downto 0);
 subtype U_Word              is UNSIGNED (15 downto 0);
 subtype U_Seventeen_Bits    is UNSIGNED (16 downto 0);
 subtype U_Eigthteen_Bits    is UNSIGNED (17 downto 0);
 subtype U_Nineteen_Bits     is UNSIGNED (18 downto 0);
 subtype U_Twenty_Bits       is UNSIGNED (19 downto 0);
 subtype U_Twenty1_Bits	     is UNSIGNED (20 downto 0);
 subtype U_Twenty2_Bits      is UNSIGNED (21 downto 0);
 subtype U_Twenty3_Bits      is UNSIGNED (22 downto 0);
 subtype U_Twenty4_Bits      is UNSIGNED (23 downto 0);
 subtype U_Twenty5_Bits      is UNSIGNED (24 downto 0);
 subtype U_Twenty6_Bits      is UNSIGNED (25 downto 0);
 subtype U_Twenty7_Bits      is UNSIGNED (26 downto 0);
 subtype U_Twenty8_Bits      is UNSIGNED (27 downto 0);
 subtype U_Twenty9_Bits      is UNSIGNED (28 downto 0);
 subtype U_Thirty_Bits       is UNSIGNED (29 downto 0);
 subtype U_Thirty1_Bits      is UNSIGNED (30 downto 0);
 subtype U_Long_Word         is UNSIGNED (31 downto 0);
 subtype U_Thirty3_Bits      is UNSIGNED (32 downto 0);
 subtype U_Thirty4_Bits      is UNSIGNED (33 downto 0);
 subtype U_Thirty5_Bits      is UNSIGNED (34 downto 0);
 subtype U_Thirty6_Bits      is UNSIGNED (35 downto 0);
 subtype U_Thirty7_Bits      is UNSIGNED (36 downto 0);
 subtype U_Thirty8_Bits      is UNSIGNED (37 downto 0);
 subtype U_Thirty9_Bits      is UNSIGNED (38 downto 0);
 subtype U_Forty_Bits       is UNSIGNED (39 downto 0);
 subtype U_Forty1_Bits      is UNSIGNED (40 downto 0);
 subtype U_Forty2_Bits      is UNSIGNED (41 downto 0);
 subtype U_Forty3_Bits      is UNSIGNED (42 downto 0);
 subtype U_Forty4_Bits      is UNSIGNED (43 downto 0);
 subtype U_Forty5_Bits      is UNSIGNED (44 downto 0);
--
 subtype S_Two_Bits          is SIGNED (1 downto 0);
 subtype S_Three_Bits        is SIGNED (2 downto 0);
 subtype S_NIBBLE            is SIGNED (3 downto 0);
 subtype S_Five_Bits         is SIGNED (4 downto 0);
 subtype S_Six_Bits          is SIGNED (5 downto 0);
 subtype S_Seven_Bits        is SIGNED (6 downto 0);
 subtype S_Byte              is SIGNED (7 downto 0);
 subtype S_Nine_Bits         is SIGNED (8 downto 0);
 subtype S_Ten_Bits          is SIGNED (9 downto 0);
 subtype S_Eleven_Bits       is SIGNED (10 downto 0);
 subtype S_Twelve_Bits       is SIGNED (11 downto 0);
 subtype S_Thirteen_Bits     is SIGNED (12 downto 0);
 subtype S_Fourteen_Bits     is SIGNED (13 downto 0);
 subtype S_Fifteen_Bits      is SIGNED (14 downto 0);
 subtype S_Word              is SIGNED (15 downto 0);
 subtype S_Seventeen_Bits    is SIGNED (16 downto 0);
 subtype S_Eigthteen_Bits    is SIGNED (17 downto 0);
 subtype S_Nineteen_Bits     is SIGNED (18 downto 0);
 subtype S_Twenty_Bits       is SIGNED (19 downto 0);
 subtype S_Twenty1_Bits	     is SIGNED (20 downto 0);
 subtype S_Twenty2_Bits      is SIGNED (21 downto 0);
 subtype S_Twenty3_Bits      is SIGNED (22 downto 0);
 subtype S_Twenty4_Bits      is SIGNED (23 downto 0);
 subtype S_Twenty5_Bits      is SIGNED (24 downto 0);
 subtype S_Twenty6_Bits      is SIGNED (25 downto 0);
 subtype S_Twenty7_Bits      is SIGNED (26 downto 0);
 subtype S_Twenty8_Bits      is SIGNED (27 downto 0);
 subtype S_Twenty9_Bits      is SIGNED (28 downto 0);
 subtype S_Thirty_Bits       is SIGNED (29 downto 0);
 subtype S_Thirty1_Bits      is SIGNED (30 downto 0);
 subtype S_Long_Word         is SIGNED (31 downto 0);
 subtype S_Thirty3_Bits      is SIGNED (32 downto 0);
 subtype S_Thirty4_Bits      is SIGNED (33 downto 0);
 subtype S_Thirty5_Bits      is SIGNED (34 downto 0);
 subtype S_Thirty6_Bits      is SIGNED (35 downto 0);
 subtype S_Thirty7_Bits      is SIGNED (36 downto 0);
 subtype S_Thirty8_Bits      is SIGNED (37 downto 0);
 subtype S_Thirty9_Bits      is SIGNED (38 downto 0);
 subtype S_Forty_Bits       is SIGNED (39 downto 0);
 subtype S_Forty1_Bits      is SIGNED (40 downto 0);
 subtype S_Forty2_Bits      is SIGNED (41 downto 0);
 subtype S_Forty3_Bits      is SIGNED (42 downto 0);
 subtype S_Forty4_Bits      is SIGNED (43 downto 0);
 subtype S_Forty5_Bits      is SIGNED (44 downto 0);
--
 
end package MATRIX_PACKAGE;

Library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY MUL_1 IS
PORT (A, B : IN UNSIGNED; Z : OUT UNSIGNED);
END ENTITY;

ARCHITECTURE BEHAVIOURAL OF MUL_1 IS
BEGIN 
        Z <= A + B;
        
END ARCHITECTURE BEHAVIOURAL;

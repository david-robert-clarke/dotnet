-- FINAL YEAR PROJECT MARK III
-- BY DAVID.R.CLARKE
-- DATE 8_12_2000
-- UPDATED ON 11_12_2000
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEe.STD_LOGIC_ARITH.ALL;
USE WORK.MATRIX_PACKAGE.ALL;
--
ENTITY MUL2 IS
PORT (A, B : IN U_TWO_BITS; Z : OUT NIBBLE);
END ENTITY MUL2;
-- 
ARCHITECTURE BEHAVIOURAL OF MUL2 IS
SIGNAL A0, B0 : ONE_BIT;
BEGIN
	Z  <= CONV_STD_LOGIC_VECTOR((A*B), 4);
	 
END ARCHITECTURE BEHAVIOURAL;

-- CREATED BY DAVID CLARKE ON 30_11_2000
-- FOR THE FINAL YEAR PROJECT
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
--
ENTITY PART_LATCH_A IS
PORT (PART_OUT : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      CLK : IN STD_LOGIC; A_LATCH_EN : IN STD_LOGIC;
      A_OUT : OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END PART_LATCH_A;
--
ARCHITECTURE STRUCTURAL OF PART_LATCH_A IS

BEGIN 

END ARCHITECTURE STRUCTURAL;

-- CREATED BY DAVID CLARKE ON 30_11_2000
-- FOR THE FINAL YEAR PROJECT
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
--
ENTITY EN_DEC IS
PORT (LATCHES_EN : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      A_LATCH_EN, B_LATCH_EN, C_LATCH_EN, D_LATCH_EN : OUT STD_lOGIC);
END ENTITY EN_DEC;

ARCHITECTURE BEHAVIOURAL OF EN_DEC IS
BEGIN
    
    SPLIT : PROCESS (LATCHES_EN) IS
    BEGIN
        IF LATCHES_EN = "11" THEN
           A_LATCH_EN <= '1'; B_LATCH_EN <= '0'; C_LATCH_EN <= '0'; 
           D_LATCH_EN <= '0';
        ELSIF LATCHES_EN = "10" THEN
           A_LATCH_EN <= '0'; B_LATCH_EN <= '1'; C_LATCH_EN <= '0'; 
           D_LATCH_EN <= '0';
        ELSIF LATCHES_EN = "01" THEN
           A_LATCH_EN <= '0'; B_LATCH_EN <= '0'; C_LATCH_EN <= '1'; 
           D_LATCH_EN <= '0';
        ELSIF LATCHES_EN = "00" THEN
           A_LATCH_EN <= '0'; B_LATCH_EN <= '0'; C_LATCH_EN <= '0'; 
           D_LATCH_EN <= '1';
        END IF;
    END PROCESS SPLIT;
    
END ARCHITECTURE BEHAVIOURAL;

-- Behavioural 32x7 ROM 
-- Final Year Project
-- By David Clarke
-- Created on 07_02_2001

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
USE WORK.MATRIX_PACKAGE.ALL;
--
entity data_store is
     port (ADDR_31, ADDR_30, ADDR_29, ADDR_28, ADDR_27, ADDR_26, ADDR_25, ADDR_24, 
           ADDR_23, ADDR_22, ADDR_21, ADDR_20, ADDR_19, ADDR_18, ADDR_17, ADDR_16, 
           ADDR_15, ADDR_14, ADDR_13, ADDR_12, ADDR_11, ADDR_10, ADDR_9, ADDR_8,
           ADDR_7, ADDR_6, ADDR_5, ADDR_4, ADDR_3, ADDR_2, ADDR_1, ADDR_0: in unsigned(1 downto 0);
           A11, A12, A13, A14, B11, B12, B13, B14,
     	   A21, A22, A23, A24, B21, B22, B23, B24,
     	   A31, A32, A33, A34, B31, B32, B33, B34,
     	   A41, A42, A43, A44, B41, B42, B43, B44  : OUT U_TWO_BITS);
end data_store;

architecture Behavioural of data_store is
    subtype ROM_BITS is U_TWO_BITS;
    type ROM_TABLE is array (3 downto 0) of ROM_BITS;
    constant ROM: ROM_TABLE := ROM_TABLE'(ROM_BITS'("11"), ROM_BITS'("10"), ROM_BITS'("01"), ROM_BITS'("00"));
                                        
begin 

-- THIS SYSTEM USES THE CONV_INTEGER FUNCTION TO CONVERT THE ADDRESS FROM A LOGIC VALUE TO AN INTEGER IN ORDER
-- TO BE USED TO ADDRESS THE REQUIRED MEMORY BITS

        A11 <= ROM(CONV_INTEGER(ADDR_31));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_31
        A12 <= ROM(CONV_INTEGER(ADDR_30));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_30
        A13 <= ROM(CONV_INTEGER(ADDR_29));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_29
        A14 <= ROM(CONV_INTEGER(ADDR_28));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_28
        A21 <= ROM(CONV_INTEGER(ADDR_27));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_27
        A22 <= ROM(CONV_INTEGER(ADDR_26));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_26
        A23 <= ROM(CONV_INTEGER(ADDR_25));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_25
        A24 <= ROM(CONV_INTEGER(ADDR_24));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_24
        A31 <= ROM(CONV_INTEGER(ADDR_23));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_23
        A32 <= ROM(CONV_INTEGER(ADDR_22));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_22
        A33 <= ROM(CONV_INTEGER(ADDR_21));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_21
        A34 <= ROM(CONV_INTEGER(ADDR_20));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_20
        A41 <= ROM(CONV_INTEGER(ADDR_19));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_19
        A42 <= ROM(CONV_INTEGER(ADDR_18));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_18
        A43 <= ROM(CONV_INTEGER(ADDR_17));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_17
        A44 <= ROM(CONV_INTEGER(ADDR_16));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_16
        B11 <= ROM(CONV_INTEGER(ADDR_15));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_15
        B12 <= ROM(CONV_INTEGER(ADDR_14));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_14
        B13 <= ROM(CONV_INTEGER(ADDR_13));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_13
        B14 <= ROM(CONV_INTEGER(ADDR_12));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_12
        B21 <= ROM(CONV_INTEGER(ADDR_11));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_11
        B22 <= ROM(CONV_INTEGER(ADDR_10));  -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_10
        B23 <= ROM(CONV_INTEGER(ADDR_9));   -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_9
        B24 <= ROM(CONV_INTEGER(ADDR_8));   -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_8
        B31 <= ROM(CONV_INTEGER(ADDR_7));   -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_7
        B32 <= ROM(CONV_INTEGER(ADDR_6));   -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_6
        B33 <= ROM(CONV_INTEGER(ADDR_5));   -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_5
        B34 <= ROM(CONV_INTEGER(ADDR_4));   -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_4
        B41 <= ROM(CONV_INTEGER(ADDR_3));   -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_3
        B42 <= ROM(CONV_INTEGER(ADDR_2));   -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_2
        B43 <= ROM(CONV_INTEGER(ADDR_1));   -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_1
        B44 <= ROM(CONV_INTEGER(ADDR_0));   -- READ FROM THE ROM USING A TWO BIT ADDRESS LINE ADDR_0
 
end Behavioural;


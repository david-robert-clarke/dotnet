-- Created by David Clarke
-- Final Year Project
-- Exploiting Parallelism in FPGA design
-- Date : 4_12_2000
Library IEEE;
Use IEEE.STD_LOGIC_1164.ALL;

ENTITY config2_latches IS
PORT (PARTITION_OUT : IN STD_LOGIC_VECTOR (15 downto 0);
      CLK, CLR      : IN STD_LOGIC;
      MUX_SEL       : IN STD_LOGIC_VECTOR (1 downto 0);
      LATCH_OUT     : OUT STD_LOGIC_VECTOR (15 downto 0));
END ENTITY config2_latches;

ARCHITECTURE Structural OF config2_latches IS

COMPONENT En_Conflict_Res_Mux2 IS
PORT (IN1, IN0 : IN STD_LOGIC; OUT1 : OUT STD_LOGIC);
END COMPONENT En_Conflict_Res_Mux2;

COMPONENT En_Conflict_Res_Mux3 IS
PORT (IN2, IN1, IN0 : IN STD_LOGIC; OUT1 : OUT STD_LOGIC);
END COMPONENT En_Conflict_Res_Mux3;

COMPONENT FDCE IS
PORT (D, CLK, CLR, CE : IN STD_LOGIC; Q : OUT STD_LOGIC);
END COMPONENT FDCE;

COMPONENT MUX_SEL3 IS
PORT (D_LATCH : IN STD_LOGIC; EXT_DATA : IN STD_LOGIC_VECTOR (1 downto 0);
      SEL : IN STD_LOGIC_VECTOR (1 downto 0); Q : OUT STD_LOGIC);
END COMPONENT MUX_SEL3;

COMPONENT MUX_SEL2 IS
PORT (D_LATCH, EXT_DATA : IN STD_LOGIC; 
      SEL : IN STD_LOGIC_VECTOR (1 downto 0); Q : OUT STD_LOGIC);
END COMPONENT MUX_SEL2;

COMPONENT Latch_En_Dec IS
PORT (INPUT : IN STD_LOGIC_VECTOR (1 downto 0) ; LATCH_EN_1, LATCH_EN_2, 
      LATCH_EN_3 : OUT STD_LOGIC);
END COMPONENT Latch_En_Dec;

SIGNAL AI, AO, BI, BO, CI, CO, DI, DO, EI, EO, FI, FO, GI, GO, HI, HO, II, IO, JI, JO, 
       KI, KO, LI, LO, MI, MO, NI, NO, OI, OO, PI, PO, EN_1, EN_2, EN_3, EN21_24, EN11_14, EN15_18 : STD_LOGIC;

BEGIN
    
    -- LOOKING AT THE SCHEMATIC CREATED IN MICROSOFT WORD, THE VHDL STRUCTURAL CODE FOLLOWS THE LAYOUT
    -- FROM THE LEFT TO THE RIGHT SIDE OF THE PAGE
    
    DEATH    : Latch_En_Dec PORT MAP (INPUT => MUX_SEL, LATCH_EN_1 => EN_1, LATCH_EN_2 => EN_2, LATCH_EN_3 => EN_3); 
    
    RES21_24 : En_Conflict_Res_Mux2 PORT MAP (IN1 => EN_2, IN0 => EN_1, OUT1 => EN21_24);
    RES15_18 : En_Conflict_Res_Mux2 PORT MAP (IN1 => EN_3, IN0 => EN_2, OUT1 => EN15_18);
    RES11_14 : En_Conflict_Res_Mux3 PORT MAP (IN2 => EN_3, IN1 => EN_2, IN0 => EN_1, OUT1 => EN11_14);
    
    DFF41 : FDCE PORT MAP (D => PARTITION_OUT(3), CLK => CLK, CLR => CLR, CE => EN_1, Q => AI);
    DFF42 : FDCE PORT MAP (D => PARTITION_OUT(2), CLK => CLK, CLR => CLR, CE => EN_1, Q => BI);
    DFF43 : FDCE PORT MAP (D => PARTITION_OUT(1), CLK => CLK, CLR => CLR, CE => EN_1, Q => CI);
    DFF44 : FDCE PORT MAP (D => PARTITION_OUT(0), CLK => CLK, CLR => CLR, CE => EN_1, Q => DI);
    
    MUXA  : MUX_SEL2 PORT MAP (D_LATCH => AI, EXT_DATA => PARTITION_OUT(7), SEL => MUX_SEL, Q => AO);
    MUXB  : MUX_SEL2 PORT MAP (D_LATCH => BI, EXT_DATA => PARTITION_OUT(6), SEL => MUX_SEL, Q => BO);
    MUXC  : MUX_SEL2 PORT MAP (D_LATCH => CI, EXT_DATA => PARTITION_OUT(5), SEL => MUX_SEL, Q => CO);
    MUXD  : MUX_SEL2 PORT MAP (D_LATCH => DI, EXT_DATA => PARTITION_OUT(4), SEL => MUX_SEL, Q => DO);
    
    DFF31 : FDCE PORT MAP (D => AO, CLK => CLK, CLR => CLR, CE => EN_1, Q => EI);
    DFF32 : FDCE PORT MAP (D => BO, CLK => CLK, CLR => CLR, CE => EN_1, Q => FI);
    DFF33 : FDCE PORT MAP (D => CO, CLK => CLK, CLR => CLR, CE => EN_1, Q => GI);
    DFF34 : FDCE PORT MAP (D => DO, CLK => CLK, CLR => CLR, CE => EN_1, Q => HI);
    
    MUXE  : MUX_SEL3 PORT MAP (D_LATCH => EI, EXT_DATA(1) => PARTITION_OUT(11), EXT_DATA(0) => PARTITION_OUT(7), 
                               SEL => MUX_SEL, Q => EO);
    MUXF  : MUX_SEL3 PORT MAP (D_LATCH => FI, EXT_DATA(1) => PARTITION_OUT(10), EXT_DATA(0) => PARTITION_OUT(6), 
                               SEL => MUX_SEL, Q => FO);
    MUXG  : MUX_SEL3 PORT MAP (D_LATCH => GI, EXT_DATA(1) => PARTITION_OUT(9),  EXT_DATA(0) => PARTITION_OUT(5), 
                               SEL => MUX_SEL, Q => GO);
    MUXH  : MUX_SEL3 PORT MAP (D_LATCH => HI, EXT_DATA(1) => PARTITION_OUT(8),  EXT_DATA(0) => PARTITION_OUT(4), 
                               SEL => MUX_SEL, Q => HO);
                               
    DFF21 : FDCE PORT MAP (D => EO, CLK => CLK, CLR => CLR, CE => EN21_24, Q => II);
    DFF22 : FDCE PORT MAP (D => FO, CLK => CLK, CLR => CLR, CE => EN21_24, Q => JI);
    DFF23 : FDCE PORT MAP (D => GO, CLK => CLK, CLR => CLR, CE => EN21_24, Q => KI);
    DFF24 : FDCE PORT MAP (D => HO, CLK => CLK, CLR => CLR, CE => EN21_24, Q => LI);
    DFF25 : FDCE PORT MAP (D => PARTITION_OUT(3), CLK => CLK, CLR => CLR, CE => EN_2, Q => MI);
    DFF26 : FDCE PORT MAP (D => PARTITION_OUT(2), CLK => CLK, CLR => CLR, CE => EN_2, Q => NI);
    DFF27 : FDCE PORT MAP (D => PARTITION_OUT(1), CLK => CLK, CLR => CLR, CE => EN_2, Q => OI);
    DFF28 : FDCE PORT MAP (D => PARTITION_OUT(0), CLK => CLK, CLR => CLR, CE => EN_2, Q => PI);
    
    MUXI  : MUX_SEL2 PORT MAP (D_LATCH => II, EXT_DATA => PARTITION_OUT(15), SEL => MUX_SEL, Q => IO);
    MUXJ  : MUX_SEL2 PORT MAP (D_LATCH => JI, EXT_DATA => PARTITION_OUT(14), SEL => MUX_SEL, Q => JO);
    MUXK  : MUX_SEL2 PORT MAP (D_LATCH => KI, EXT_DATA => PARTITION_OUT(13), SEL => MUX_SEL, Q => KO);
    MUXL  : MUX_SEL2 PORT MAP (D_LATCH => LI, EXT_DATA => PARTITION_OUT(12), SEL => MUX_SEL, Q => LO);
    MUXM  : MUX_SEL2 PORT MAP (D_LATCH => MI, EXT_DATA => PARTITION_OUT(11), SEL => MUX_SEL, Q => MO);
    MUXN  : MUX_SEL2 PORT MAP (D_LATCH => NI, EXT_DATA => PARTITION_OUT(10), SEL => MUX_SEL, Q => NO);
    MUXO  : MUX_SEL2 PORT MAP (D_LATCH => OI, EXT_DATA => PARTITION_OUT(9),  SEL => MUX_SEL, Q => OO);
    MUXP  : MUX_SEL2 PORT MAP (D_LATCH => PI, EXT_DATA => PARTITION_OUT(8),  SEL => MUX_SEL, Q => PO);
    
    DFF11 : FDCE PORT MAP (D => IO, CLK => CLK, CLR => CLR, CE => EN11_14, Q => LATCH_OUT(15));
    DFF12 : FDCE PORT MAP (D => JO, CLK => CLK, CLR => CLR, CE => EN11_14, Q => LATCH_OUT(14));
    DFF13 : FDCE PORT MAP (D => KO, CLK => CLK, CLR => CLR, CE => EN11_14, Q => LATCH_OUT(13));
    DFF14 : FDCE PORT MAP (D => LO, CLK => CLK, CLR => CLR, CE => EN11_14, Q => LATCH_OUT(12));
    DFF15 : FDCE PORT MAP (D => MO, CLK => CLK, CLR => CLR, CE => EN15_18, Q => LATCH_OUT(11));
    DFF16 : FDCE PORT MAP (D => NO, CLK => CLK, CLR => CLR, CE => EN15_18, Q => LATCH_OUT(10));
    DFF17 : FDCE PORT MAP (D => OO, CLK => CLK, CLR => CLR, CE => EN15_18, Q => LATCH_OUT(9));
    DFF18 : FDCE PORT MAP (D => PO, CLK => CLK, CLR => CLR, CE => EN15_18, Q => LATCH_OUT(8));
    DFF19 : FDCE PORT MAP (D => PARTITION_OUT(7), CLK => CLK, CLR => CLR, CE => EN_3, Q => LATCH_OUT(7));
    DFF1A : FDCE PORT MAP (D => PARTITION_OUT(6), CLK => CLK, CLR => CLR, CE => EN_3, Q => LATCH_OUT(6));
    DFF1B : FDCE PORT MAP (D => PARTITION_OUT(5), CLK => CLK, CLR => CLR, CE => EN_3, Q => LATCH_OUT(5));
    DFF1C : FDCE PORT MAP (D => PARTITION_OUT(4), CLK => CLK, CLR => CLR, CE => EN_3, Q => LATCH_OUT(4));
    DFF1D : FDCE PORT MAP (D => PARTITION_OUT(3), CLK => CLK, CLR => CLR, CE => EN_3, Q => LATCH_OUT(3));
    DFF1E : FDCE PORT MAP (D => PARTITION_OUT(2), CLK => CLK, CLR => CLR, CE => EN_3, Q => LATCH_OUT(2));
    DFF1F : FDCE PORT MAP (D => PARTITION_OUT(1), CLK => CLK, CLR => CLR, CE => EN_3, Q => LATCH_OUT(1));
    DFF1G : FDCE PORT MAP (D => PARTITION_OUT(0), CLK => CLK, CLR => CLR, CE => EN_3, Q => LATCH_OUT(0));
                              
END ARCHITECTURE Structural;

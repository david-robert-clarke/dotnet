-- Final Year Project
-- By David.R.Clarke
-- Created 20_12_2000
Library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE WORK.MATRIX_PACKAGE.ALL;
ENTITY SYSTEMS_123 IS
PORT (signal RESET, CLK : IN ONE_BIT;
      A0B0_A1B2_CONFIG_3, A0B0_A1B2_CONFIG_2, A0B0_A1B2_CONFIG_1,
      A0B1_A1B3_CONFIG_3, A0B1_A1B3_CONFIG_2, A0B1_A1B3_CONFIG_1,
      A2B0_A3B2_CONFIG_3, A2B0_A3B2_CONFIG_2, A2B0_A3B2_CONFIG_1,
      A2B1_A3B3_CONFIG_3, A2B1_A3B3_CONFIG_2, A2B1_A3B3_CONFIG_1 : OUT FIVE_BITS);
END ENTITY SYSTEMS_123;
--
ARCHITECTURE STRUCTURAL OF SYSTEMS_123 IS

component STARTUP
  port (GSR: in std_logic);
end component;

COMPONENT SYSTEM_3 is
     Port (CLK, RESET : IN ONE_BIT;
           A0B0_A1B2, A0B1_A1B3, A2B0_A3B2, A2B1_A3B3 : OUT FIVE_BITS);
End COMPONENT SYSTEM_3;

COMPONENT SYSTEM_2 is
     Port (CLK, RESET : IN ONE_BIT;
           A0B0_A1B2, A0B1_A1B3, A2B0_A3B2, A2B1_A3B3 : OUT FIVE_BITS);
End COMPONENT SYSTEM_2;

COMPONENT SYSTEM is
     Port (CLK, RESET : IN ONE_BIT;
           A0B0_A1B2, A0B1_A1B3, A2B0_A3B2, A2B1_A3B3 : OUT FIVE_BITS);
End COMPONENT SYSTEM;

SIGNAL GSR_NET : ONE_BIT;

BEGIN

U1: STARTUP  port map (GSR=>RESET);

CONFIG_3 : SYSTEM_3 PORT MAP (CLK => CLK, RESET => RESET, A0B0_A1B2 => A0B0_A1B2_CONFIG_3, A0B1_A1B3 => A0B1_A1B3_CONFIG_3, 
                              A2B0_A3B2 => A2B0_A3B2_CONFIG_3, A2B1_A3B3 => A2B1_A3B3_CONFIG_3);
CONFIG_2 : SYSTEM_2 PORT MAP (CLK => CLK, RESET => RESET, A0B0_A1B2 => A0B0_A1B2_CONFIG_2, A0B1_A1B3 => A0B1_A1B3_CONFIG_2, 
                              A2B0_A3B2 => A2B0_A3B2_CONFIG_2, A2B1_A3B3 => A2B1_A3B3_CONFIG_2);
CONFIG_1 : SYSTEM   PORT MAP (CLK => CLK, RESET => RESET, A0B0_A1B2 => A0B0_A1B2_CONFIG_1, A0B1_A1B3 => A0B1_A1B3_CONFIG_1, 
                              A2B0_A3B2 => A2B0_A3B2_CONFIG_1, A2B1_A3B3 => A2B1_A3B3_CONFIG_1);
END ARCHITECTURE STRUCTURAL;










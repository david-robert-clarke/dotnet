-- Created by David Clarke for the RS232 assignment
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

Entity AND4B2 IS
Port (a, b, c, d : IN std_logic; z : OUT std_logic);
End Entity AND4B2;

Architecture Behavioural OF AND4B2 IS
Begin
   z <= a AND b AND (NOT c) AND (NOT d);
End Architecture Behavioural;

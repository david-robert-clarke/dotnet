-- Final Year Project
-- By David Clarke
-- Created: 16_12_2000
Entity MEM_EL IS
PORT
End Entity MEM_EL;
--
Architecture Behavioural of MEM_EL is
Begin
End Architecture Behavioural;

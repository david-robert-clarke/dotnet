-- CREATED BY DAVID CLARKE ON 30_11_2000
-- FOR THE FINAL YEAR PROJECT
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
--
ENTITY PART_LATCH_D IS
PORT (PART_OUT : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      CLK : IN STD_LOGIC; D_LATCH_EN : IN STD_LOGIC;
      D_OUT : OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END PART_LATCH_D;
--
ARCHITECTURE STRUCTURAL OF PART_LATCH_D IS

BEGIN 

END ARCHITECTURE STRUCTURAL;

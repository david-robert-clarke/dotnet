-- Test material
Library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE WORK.MATRIX_PACKAGE.ALL;
--
ENTITY ADDER_4_BIT IS
PORT (A, B : IN U_NIBBLE; Z : OUT U_NIBBLE);
END ENTITY ADDER_4_BIT;

ARCHITECTURE BEHAVIOURAL OF ADDER_4_BIT IS
BEGIN
	Z <= A + B;
END ARCHITECTURE BEHAVIOURAL; 

-- Final Year Project MarkIII
-- Created by David.R.Clarke
-- Date: 9_12_2000
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
--
ENTITY ADD4 IS
PORT (A, B : IN STD_LOGIC_VECTOR (3 downto 0);
      S : OUT STD_LOGIC_VECTOR (3 downto 0); COUT : OUT STD_LOGIC);
END ENTITY ADD4;
--
ARCHITECTURE STRUCTURAL OF ADD4 IS

COMPONENT FULL_ADDER IS
PORT (A, B, C_IN : IN std_logic; 
      SUM, C_OUT : OUT std_logic);
END COMPONENT FULL_ADDER; 

COMPONENT FULL_ADDERIN IS
PORT (A, B : IN std_logic; 
      SUM, C_OUT : OUT std_logic);
END COMPONENT FULL_ADDERIN; 

SIGNAL COCI1_2, COCI2_3, COCI3_4 : STD_LOGIC; 

BEGIN

ADDERN01 : FULL_ADDERIN PORT MAP (A => A(0), B => B(0), SUM => S(0), C_OUT => COCI1_2);
ADDERN02 : FULL_ADDER   PORT MAP (A => A(1), B => B(1), C_IN => COCI1_2, SUM => S(1), C_OUT => COCI2_3);
ADDERN03 : FULL_ADDER   PORT MAP (A => A(2), B => B(2), C_IN => COCI2_3, SUM => S(2), C_OUT => COCI3_4);
ADDERN04 : FULL_ADDER   PORT MAP (A => A(3), B => B(3), C_IN => COCI3_4, SUM => S(3), C_OUT => COUT);

END ARCHITECTURE STRUCTURAL;

-- Final Year Project
-- By David.R.Clarke
-- Created 14_12_2000
-- Updated 20_12_2000
Library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE WORK.MATRIX_PACKAGE.ALL;
--
Entity SYSTEM_2 is
     Port (CLK, RESET : IN ONE_BIT;
           A0B0_A1B2, A0B1_A1B3, A2B0_A3B2, A2B1_A3B3 : OUT FIVE_BITS);
End Entity SYSTEM_2;

Architecture STRUCTURAL of SYSTEM_2 is
-- Component Declarations

--Component STARTUP
--Port (GSR: in std_logic);
--End Component;

Component DSP_CONFIG_2 IS
Port (C, R : IN ONE_BIT;
      MAT_A_D_IN_3, MAT_A_D_IN_2, MAT_A_D_IN_1, MAT_A_D_IN_0,  
      MAT_B_D_IN_3, MAT_B_D_IN_2, MAT_B_D_IN_1, MAT_B_D_IN_0 : IN U_TWO_BITS;
      SEL : IN ONE_BIT; A0B0_A1B2, A0B1_A1B3, A2B0_A3B2, A2B1_A3B3 : OUT FIVE_BITS);
End Component DSP_CONFIG_2;    

Component data_store is
Port (ADDR: in INTEGER range 1 downto 0;
      DATA: out U_WORD);
End Component data_store;

Component ASM_CONFIG_2 IS
PORT (CLK, RESET      : IN ONE_BIT; 
      DATA_SELECT     : OUT INTEGER range 1 downto 0;
      MEM_SEL_OUT     : OUT ONE_BIT);
End Component ASM_CONFIG_2;

Signal Elem_DBUS        : U_WORD;
Signal Mem_SelBus       : ONE_BIT;
Signal Data_SelBus      : INTEGER range 1 downto 0;
-- SIGNAL GSR_NET          : ONE_BIT;
Begin
-- Component Instantiations

-- U1: STARTUP  port map (GSR=>RESET);

DSP_2 : DSP_CONFIG_2          PORT MAP (C => CLK, R => RESET,
					MAT_A_D_IN_3 => Elem_DBUS(15 downto 14), MAT_B_D_IN_3 => Elem_DBUS(13 downto 12),
                                        MAT_A_D_IN_2 => Elem_DBUS(11 downto 10), MAT_B_D_IN_2 => Elem_DBUS(9 downto 8),
                                        MAT_A_D_IN_1 => Elem_DBUS(7 downto 6),   MAT_B_D_IN_1 => Elem_DBUS(5 downto 4),
                                        MAT_A_D_IN_0 => Elem_DBUS(3 downto 2),   MAT_B_D_IN_0 => Elem_DBUS(1 downto 0),
                                        SEL => Mem_SelBus, A0B0_A1B2 => A0B0_A1B2 , A0B1_A1B3 => A0B1_A1B3, 
                                        A2B0_A3B2 => A2B0_A3B2, A2B1_A3B3 => A2B1_A3B3);

Data_Store_2A  : Data_Store   PORT MAP (ADDR => Data_SelBus, DATA => Elem_DBUS);

Asm_Config_2_A : Asm_Config_2 PORT MAP (CLK => CLK, RESET => RESET, DATA_SELECT => Data_SelBus, MEM_SEL_OUT => Mem_SelBus);

End Architecture STRUCTURAL;




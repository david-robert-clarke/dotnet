-- Final Year Project
-- By David Clarke
-- Created 12_12_2000
-- Updated 14_12_2000
Library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE WORK.MATRIX_PACKAGE.ALL; -- USING MY NEW PACKAGE
--
ENTITY ASM_CONFIG_1 IS
PORT (CLK, RESET      : IN ONE_BIT; 
      DATA_SELECT     : OUT INTEGER range 3 downto 0;
      MEM_SEL_OUT     : OUT TWO_BITS);
END ENTITY ASM_CONFIG_1;
--
ARCHITECTURE STATE_MACHINE OF ASM_CONFIG_1 IS

signal CURRENT_STATE, NEXT_STATE : STATE_TYPE;

BEGIN
    next_state_logic: PROCESS (current_state) IS
         Begin   
              CASE current_state IS           
                   WHEN S0 => next_state <= S1;
                   WHEN S1 => next_state <= S2;
                   WHEN S2 => next_state <= S3;
                   WHEN S3 => next_state <= S3;
              END CASE;
         End Process next_state_logic;
        
    state_update : PROCESS (next_state, RESET, CLK) IS
         Begin
              IF rising_edge(clk) THEN
                 IF RESET = '1' THEN current_state <= S0;
                 ELSE current_state <= next_state;
                 END IF;
              END IF;
         End PROCESS state_update;
         
   output_logic : PROCESS (current_state)
        Begin
             CASE current_state IS
                  WHEN S0 =>    Data_Select <= 3; 
                  		MEM_SEL_OUT <= "11";
                  
                  WHEN S1 =>    Data_Select <= 2;
                  	        MEM_SEL_OUT <= "10";
                  
                  WHEN S2 =>	Data_Select <= 1;
                  		MEM_SEL_OUT <= "01";
                  			
                  WHEN S3 =>	Data_Select <= 0;
                  		MEM_SEL_OUT <= "00";     
             END CASE;
        END PROCESS output_logic;     
                   
END ARCHITECTURE STATE_MACHINE;
    

-- Final Year Project
-- By David Clarke
-- Created 31_01_2001
-- Updated 1_02_2001
Library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE WORK.MATRIX_PACKAGE.ALL;
--
ENTITY Answer_Store IS
PORT (EN, CLK, RESET : IN ONE_BIT; 
      INPUT : IN  UNSIGNED (95 downto 0);
      ANSWER: OUT UNSIGNED (95 downto 0));
END ENTITY Answer_Store;

ARCHITECTURE BEHAVIOURAL OF Answer_Store IS

COMPONENT STARTUP
 port (GSR : IN STD_LOGIC);
END COMPONENT STARTUP;

BEGIN

GLOBAL : STARTUP PORT MAP (GSR => RESET);

	PROCESS (INPUT, CLK, RESET, EN)
	BEGIN
	
	    IF reset = '1' THEN
	       ANSWER <= X"000000000000000000000000"; 
	    ELSE
	        IF rising_edge(CLK) THEN
	            CASE EN IS
	            WHEN '1' =>
	                ANSWER(95 downto 90) <= INPUT (95 downto 90);
	                ANSWER(89 downto 84) <= INPUT (89 downto 84);
	                ANSWER(83 downto 78) <= INPUT (83 downto 78);
	                ANSWER(77 downto 72) <= INPUT (77 downto 72);
	                ANSWER(71 downto 66) <= INPUT (71 downto 66);
	                ANSWER(65 downto 60) <= INPUT (65 downto 60);
	                ANSWER(59 downto 54) <= INPUT (59 downto 54);
	                ANSWER(53 downto 48) <= INPUT (53 downto 48);
	                ANSWER(47 downto 42) <= INPUT (47 downto 42);
	                ANSWER(41 downto 36) <= INPUT (41 downto 36);
	                ANSWER(35 downto 30) <= INPUT (35 downto 30);
	                ANSWER(29 downto 24) <= INPUT (29 downto 24);
	                ANSWER(23 downto 18) <= INPUT (23 downto 18);
	                ANSWER(17 downto 12) <= INPUT (17 downto 12);
	                ANSWER(11 downto 6)  <= INPUT (11 downto 6);
	                ANSWER(5 downto 0)   <= INPUT (5 downto 0);
	            WHEN OTHERS =>
	                 NULL;
	            END CASE;
	       END IF;
	    END IF;
	END PROCESS;
	
END ARCHITECTURE BEHAVIOURAL;
	        
	        

-- FINAL YEAR PROJECT MARK III
-- BY DAVID.R.CLARKE
-- DATE 8_12_2000
-- UPDATED ON 11_12_2000
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEe.STD_LOGIC_ARITH.ALL;
--
ENTITY MUL2 IS
PORT (A, B : UNSIGNED (1 downto 0); Z : OUT STD_LOGIC_VECTOR (3 downto 0));
END ENTITY MUL2;
-- 
ARCHITECTURE BEHAVIOURAL OF MUL2 IS
SIGNAL A0, B0 : STD_LOGIC;
BEGIN
	-- A0 <= CONV_UNSIGNED(A,  1) ;
	-- B0 <= CONV_UNSIGNED(B,  1) ;
	Z  <= CONV_STD_LOGIC_VECTOR((A*B), 4);
	 
END ARCHITECTURE BEHAVIOURAL;

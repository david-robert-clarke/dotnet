-- Created by David Clarke
-- Final Year Project
-- Exploiting Parallelism in FPGA design
-- Date : 5_12_2000
Library IEEE;
Use IEEE.STD_LOGIC_1164.ALL;

ENTITY PART_SYNC IS
PORT (CLK, CLR : IN STD_LOGIC;
      MAT_IN : IN STD_LOGIC_VECTOR (3 downto 0);
      PARTITION_OUT : OUT STD_LOGIC_VECTOR (15 downto 0));
END ENTITY PART_SYNC;
--
ARCHITECTURE STRUCTURAL OF PART_SYNC IS

COMPONENT PART_DEC IS
PORT (INPUT : IN STD_LOGIC_VECTOR (3 downto 0);
      OUTPUT : OUT STD_LOGIC_VECTOR (15 downto 0));
END COMPONENT PART_DEC;

COMPONENT PART_LATCHES IS
PORT (CLK, CLR : IN STD_LOGIC;
      A, B, C, D : IN STD_LOGIC_VECTOR (3 downto 0); 
      Z : OUT STD_LOGIC_VECTOR (15 downto 0));
END COMPONENT PART_LATCHES;

SIGNAL PART_IN_SIG : STD_LOGIC_VECTOR (15 downto 0); 

BEGIN

PART_DEC1     : PART_DEC     PORT MAP (INPUT => MAT_IN, OUTPUT => PART_IN_SIG);
PART_LATCHES1 : PART_LATCHES PORT MAP (CLK => CLK, CLR => CLR, A => PART_IN_SIG(15 DOWNTO 12),
                                       B => PART_IN_SIG(11 DOWNTO 8), C => PART_IN_SIG(7 DOWNTO 4),
                                       D => PART_IN_SIG(3 DOWNTO 0), Z => PARTITION_OUT);
END ARCHITECTURE STRUCTURAL;

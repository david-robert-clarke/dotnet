-- Final Year Project Messaround
-- Created by David Clarke
library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
--						 
ENTITY DECODER IS
	PORT (SEL : IN STD_LOGIC_VECTOR (3 downto 0); 
	      DATA: OUT UNSIGNED (63 downto 0));
END ENTITY DECODER;

ARCHITECTURE BEHAVIOURAL OF DECODER IS

BEGIN
	GET_OUTPUT : PROCESS (SEL)
	BEGIN  
		CASE SEL IS
			WHEN "0000" 	=> DATA <= X"1111111100000001";
			WHEN "0001"	=> DATA <= X"0111111100000001";
			WHEN "0010"	=> DATA <= X"0011111100000001";
			WHEN "0011"	=> DATA <= X"0001111100000001";
			WHEN "0100"	=> DATA <= X"0000111100000001";
			WHEN "0101"	=> DATA <= X"0000011100000001";
			WHEN "0110"	=> DATA <= X"0000001100000001";
			WHEN "0111"	=> DATA <= X"0000000100000001";	
			WHEN "1000"	=> DATA <= X"0000000000000001";
			WHEN "1001"	=> DATA <= X"1111111100000000";
			WHEN "1010"	=> DATA <= X"1111111100000010";
			WHEN "1011"	=> DATA <= X"1111111100000110";
			WHEN "1100"	=> DATA <= X"1111111100001110";
			WHEN "1101"	=> DATA <= X"1111111100011110";
			WHEN "1110" 	=> DATA <= X"1111111100111110";
			WHEN OTHERS 	=> DATA <= X"1111111101111110";	   
		END CASE;
	END PROCESS GET_OUTPUT;
		
END BEHAVIOURAL;
